../.././../test/execute_tb.sv
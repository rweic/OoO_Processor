../../src/verilog/PARAM.vh
# 
# LEF OUT API 
# User Name : gbeatty3 
# Date : Mon Jun  5 00:39:42 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

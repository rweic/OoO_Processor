module issue ();
    input clk, reset;

    // Read ready operands


    // For not ready operands, rename it 




endmodule
/* Decode Module
 * pre-assign resource, rename reg to solve data dependencies
 */
module decode ();
    input clk_i, reset_i;

    // decoder dec0 ();

endmodule
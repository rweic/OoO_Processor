../../src/verilog/fsm.sv
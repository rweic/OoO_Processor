module issue ();
    input clk_i, reset_i;
    input [31:0] pc_i;
    // Should include the data that load/ store needs, or the original inst
    input [31:0] inst_i;

    // Read ready operands


    // For not ready operands, rename it 




endmodule
module decode ();
    input clk_i, reset_i;

    // decoder dec0 ();

endmodule
/* Register Rename
 * The module was supposed to solve the name dependencies
 */

module rename ();


endmodule
# 
# LEF OUT API 
# User Name : gbeatty3 
# Date : Tue May 16 23:07:53 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

# 
# LEF OUT API 
# User Name : gbeatty3 
# Date : Wed May 17 00:15:02 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

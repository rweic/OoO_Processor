../../../verilog/PARAM.vh
module muldiv_tb ();

endmodule
module fetch ();
endmodule
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO dmem
   CLASS BLOCK ;
   SIZE 235.34 BY 144.62 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.0 0.0 42.14 0.42 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  45.08 0.0 45.22 0.42 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.88 0.0 48.02 0.42 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.68 0.0 50.82 0.42 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.48 0.0 53.62 0.42 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.56 0.0 56.7 0.42 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.36 0.0 59.5 0.42 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  62.16 0.0 62.3 0.42 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.24 0.0 65.38 0.42 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  68.04 0.0 68.18 0.42 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.84 0.0 70.98 0.42 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.64 0.0 73.78 0.42 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.44 0.0 76.58 0.42 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  79.24 0.0 79.38 0.42 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.32 0.0 82.46 0.42 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  85.12 0.0 85.26 0.42 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.92 0.0 88.06 0.42 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  91.0 0.0 91.14 0.42 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.8 0.0 93.94 0.42 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.32 0.0 96.46 0.42 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.4 0.0 99.54 0.42 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  102.2 0.0 102.34 0.42 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  105.0 0.0 105.14 0.42 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.08 0.0 108.22 0.42 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.6 0.0 110.74 0.42 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.68 0.0 113.82 0.42 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.76 0.0 116.9 0.42 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.28 0.0 119.42 0.42 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  122.08 0.0 122.22 0.42 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  125.16 0.0 125.3 0.42 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  127.96 0.0 128.1 0.42 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.04 0.0 131.18 0.42 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  24.92 0.0 25.06 0.42 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  28.0 0.0 28.14 0.42 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 50.96 0.42 51.1 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 54.04 0.42 54.18 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 56.28 0.42 56.42 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 58.8 0.42 58.94 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 61.04 0.42 61.18 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 63.56 0.42 63.7 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  207.2 144.2 207.34 144.62 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  204.4 144.2 204.54 144.62 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.92 25.2 235.34 25.34 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.92 22.4 235.34 22.54 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.92 19.88 235.34 20.02 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  216.72 0.0 216.86 0.42 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  215.6 0.0 215.74 0.42 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  215.88 0.0 216.02 0.42 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 6.44 0.42 6.58 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  234.92 138.6 235.34 138.74 ;
      END
   END csb1
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.8 0.0 9.94 0.42 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  226.24 144.2 226.38 144.62 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  30.52 0.0 30.66 0.42 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.6 0.0 33.74 0.42 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.4 0.0 36.54 0.42 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  39.2 0.0 39.34 0.42 ;
      END
   END wmask0[3]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  42.56 144.2 42.7 144.62 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.04 144.2 47.18 144.62 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  51.52 144.2 51.66 144.62 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.28 144.2 56.42 144.62 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.04 144.2 61.18 144.62 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  65.8 144.2 65.94 144.62 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.28 144.2 70.42 144.62 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  75.04 144.2 75.18 144.62 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  80.08 144.2 80.22 144.62 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.84 144.2 84.98 144.62 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  89.6 144.2 89.74 144.62 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.8 144.2 93.94 144.62 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  98.84 144.2 98.98 144.62 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  103.32 144.2 103.46 144.62 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  108.36 144.2 108.5 144.62 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  112.84 144.2 112.98 144.62 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  117.32 144.2 117.46 144.62 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  122.36 144.2 122.5 144.62 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  126.84 144.2 126.98 144.62 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  131.6 144.2 131.74 144.62 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  136.36 144.2 136.5 144.62 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  141.12 144.2 141.26 144.62 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  145.88 144.2 146.02 144.62 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  150.64 144.2 150.78 144.62 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  155.12 144.2 155.26 144.62 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  159.6 144.2 159.74 144.62 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  164.64 144.2 164.78 144.62 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  169.4 144.2 169.54 144.62 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  173.88 144.2 174.02 144.62 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  178.64 144.2 178.78 144.62 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  183.12 144.2 183.26 144.62 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  187.88 144.2 188.02 144.62 ;
      END
   END dout1[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 143.22 ;
         LAYER metal3 ;
         RECT  1.4 142.52 233.94 143.22 ;
         LAYER metal3 ;
         RECT  1.4 1.4 233.94 2.1 ;
         LAYER metal4 ;
         RECT  233.24 1.4 233.94 143.22 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 0.0 235.34 0.7 ;
         LAYER metal3 ;
         RECT  0.0 143.92 235.34 144.62 ;
         LAYER metal4 ;
         RECT  234.64 0.0 235.34 144.62 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 144.62 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 235.2 144.48 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 235.2 144.48 ;
   LAYER  metal3 ;
      RECT  0.56 50.82 235.2 51.24 ;
      RECT  0.14 51.24 0.56 53.9 ;
      RECT  0.14 54.32 0.56 56.14 ;
      RECT  0.14 56.56 0.56 58.66 ;
      RECT  0.14 59.08 0.56 60.9 ;
      RECT  0.14 61.32 0.56 63.42 ;
      RECT  0.56 25.06 234.78 25.48 ;
      RECT  0.56 25.48 234.78 50.82 ;
      RECT  234.78 25.48 235.2 50.82 ;
      RECT  234.78 22.68 235.2 25.06 ;
      RECT  234.78 20.16 235.2 22.26 ;
      RECT  0.14 6.72 0.56 50.82 ;
      RECT  0.56 51.24 234.78 138.46 ;
      RECT  0.56 138.46 234.78 138.88 ;
      RECT  234.78 51.24 235.2 138.46 ;
      RECT  0.56 138.88 1.26 142.38 ;
      RECT  0.56 142.38 1.26 143.36 ;
      RECT  1.26 138.88 234.08 142.38 ;
      RECT  234.08 138.88 234.78 142.38 ;
      RECT  234.08 142.38 234.78 143.36 ;
      RECT  0.56 1.26 1.26 2.24 ;
      RECT  0.56 2.24 1.26 25.06 ;
      RECT  1.26 2.24 234.08 25.06 ;
      RECT  234.08 1.26 234.78 2.24 ;
      RECT  234.08 2.24 234.78 25.06 ;
      RECT  234.78 0.84 235.2 19.74 ;
      RECT  0.14 0.84 0.56 6.3 ;
      RECT  0.56 0.84 1.26 1.26 ;
      RECT  1.26 0.84 234.08 1.26 ;
      RECT  234.08 0.84 234.78 1.26 ;
      RECT  0.14 63.84 0.56 143.78 ;
      RECT  234.78 138.88 235.2 143.78 ;
      RECT  0.56 143.36 1.26 143.78 ;
      RECT  1.26 143.36 234.08 143.78 ;
      RECT  234.08 143.36 234.78 143.78 ;
   LAYER  metal4 ;
      RECT  42.42 0.14 44.8 0.7 ;
      RECT  45.5 0.14 47.6 0.7 ;
      RECT  48.3 0.14 50.4 0.7 ;
      RECT  51.1 0.14 53.2 0.7 ;
      RECT  53.9 0.14 56.28 0.7 ;
      RECT  56.98 0.14 59.08 0.7 ;
      RECT  59.78 0.14 61.88 0.7 ;
      RECT  62.58 0.14 64.96 0.7 ;
      RECT  65.66 0.14 67.76 0.7 ;
      RECT  68.46 0.14 70.56 0.7 ;
      RECT  71.26 0.14 73.36 0.7 ;
      RECT  74.06 0.14 76.16 0.7 ;
      RECT  76.86 0.14 78.96 0.7 ;
      RECT  79.66 0.14 82.04 0.7 ;
      RECT  82.74 0.14 84.84 0.7 ;
      RECT  85.54 0.14 87.64 0.7 ;
      RECT  88.34 0.14 90.72 0.7 ;
      RECT  91.42 0.14 93.52 0.7 ;
      RECT  94.22 0.14 96.04 0.7 ;
      RECT  96.74 0.14 99.12 0.7 ;
      RECT  99.82 0.14 101.92 0.7 ;
      RECT  102.62 0.14 104.72 0.7 ;
      RECT  105.42 0.14 107.8 0.7 ;
      RECT  108.5 0.14 110.32 0.7 ;
      RECT  111.02 0.14 113.4 0.7 ;
      RECT  114.1 0.14 116.48 0.7 ;
      RECT  117.18 0.14 119.0 0.7 ;
      RECT  119.7 0.14 121.8 0.7 ;
      RECT  122.5 0.14 124.88 0.7 ;
      RECT  125.58 0.14 127.68 0.7 ;
      RECT  128.38 0.14 130.76 0.7 ;
      RECT  25.34 0.14 27.72 0.7 ;
      RECT  42.42 0.7 206.92 143.92 ;
      RECT  206.92 0.7 207.62 143.92 ;
      RECT  204.82 143.92 206.92 144.48 ;
      RECT  131.46 0.14 215.32 0.7 ;
      RECT  216.3 0.14 216.44 0.7 ;
      RECT  10.22 0.14 24.64 0.7 ;
      RECT  207.62 143.92 225.96 144.48 ;
      RECT  28.42 0.14 30.24 0.7 ;
      RECT  30.94 0.14 33.32 0.7 ;
      RECT  34.02 0.14 36.12 0.7 ;
      RECT  36.82 0.14 38.92 0.7 ;
      RECT  39.62 0.14 41.72 0.7 ;
      RECT  41.72 0.7 42.28 143.92 ;
      RECT  41.72 143.92 42.28 144.48 ;
      RECT  42.28 0.7 42.42 143.92 ;
      RECT  42.98 143.92 46.76 144.48 ;
      RECT  47.46 143.92 51.24 144.48 ;
      RECT  51.94 143.92 56.0 144.48 ;
      RECT  56.7 143.92 60.76 144.48 ;
      RECT  61.46 143.92 65.52 144.48 ;
      RECT  66.22 143.92 70.0 144.48 ;
      RECT  70.7 143.92 74.76 144.48 ;
      RECT  75.46 143.92 79.8 144.48 ;
      RECT  80.5 143.92 84.56 144.48 ;
      RECT  85.26 143.92 89.32 144.48 ;
      RECT  90.02 143.92 93.52 144.48 ;
      RECT  94.22 143.92 98.56 144.48 ;
      RECT  99.26 143.92 103.04 144.48 ;
      RECT  103.74 143.92 108.08 144.48 ;
      RECT  108.78 143.92 112.56 144.48 ;
      RECT  113.26 143.92 117.04 144.48 ;
      RECT  117.74 143.92 122.08 144.48 ;
      RECT  122.78 143.92 126.56 144.48 ;
      RECT  127.26 143.92 131.32 144.48 ;
      RECT  132.02 143.92 136.08 144.48 ;
      RECT  136.78 143.92 140.84 144.48 ;
      RECT  141.54 143.92 145.6 144.48 ;
      RECT  146.3 143.92 150.36 144.48 ;
      RECT  151.06 143.92 154.84 144.48 ;
      RECT  155.54 143.92 159.32 144.48 ;
      RECT  160.02 143.92 164.36 144.48 ;
      RECT  165.06 143.92 169.12 144.48 ;
      RECT  169.82 143.92 173.6 144.48 ;
      RECT  174.3 143.92 178.36 144.48 ;
      RECT  179.06 143.92 182.84 144.48 ;
      RECT  183.54 143.92 187.6 144.48 ;
      RECT  188.3 143.92 204.12 144.48 ;
      RECT  1.12 0.7 2.38 1.12 ;
      RECT  1.12 143.5 2.38 144.48 ;
      RECT  2.38 0.7 41.72 1.12 ;
      RECT  2.38 1.12 41.72 143.5 ;
      RECT  2.38 143.5 41.72 144.48 ;
      RECT  207.62 0.7 232.96 1.12 ;
      RECT  207.62 1.12 232.96 143.5 ;
      RECT  207.62 143.5 232.96 143.92 ;
      RECT  232.96 0.7 234.22 1.12 ;
      RECT  232.96 143.5 234.22 143.92 ;
      RECT  217.14 0.14 234.36 0.7 ;
      RECT  226.66 143.92 234.36 144.48 ;
      RECT  234.22 0.7 234.36 1.12 ;
      RECT  234.22 1.12 234.36 143.5 ;
      RECT  234.22 143.5 234.36 143.92 ;
      RECT  0.98 0.14 9.52 0.7 ;
      RECT  0.98 0.7 1.12 1.12 ;
      RECT  0.98 1.12 1.12 143.5 ;
      RECT  0.98 143.5 1.12 144.48 ;
   END
END    dmem
END    LIBRARY

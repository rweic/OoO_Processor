module rename ();


endmodule
../../src/verilog/execute_tb.sv
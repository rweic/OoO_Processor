# 
# LEF OUT API 
# User Name : gbeatty3 
# Date : Fri May 26 19:19:14 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

# 
# LEF OUT API 
# User Name : gbeatty3 
# Date : Sun Jun  4 22:53:32 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

# 
# LEF OUT API 
# User Name : anshjsj 
# Date : Tue May  9 16:59:48 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

../../src/verilog/tb.sv
../../../test/regfile_tb.sv
../../src/verilog/toplevel_tb.sv
../../src/verilog/ram_test.sv
# 
# LEF OUT API 
# User Name : anshjsj 
# Date : Sat Apr  8 22:41:23 2023
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
END LIBRARY

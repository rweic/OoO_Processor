module decode ();
    input clk_i, reset_i;

    // module decoder ();

endmodule
../../src/verilog/alu_tb.sv
module muldiv();

endmodule
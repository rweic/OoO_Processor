../../../test/alu_tb.sv
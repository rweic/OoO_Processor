/* Mul/div Module
 * MUL lower 32 bits
 * MULH/ MULHU/ MULHSU upper 32 bits (signed×signed, unsigned×unsigned, signed×unsigned)
 * Booth Wallace Dadda Array multiplexer?
 *
 * DIV/DIVU division round towards zero
 * REM/REMU remainder (REM has the same sign as the div result)
 */
module muldiv();
    input clk_i, reset_i;
    input [31:0] pc_i;
    // Should include the data that load/ store needs, or the original inst
    input [31:0] inst_i;
    // Value of registers should be known by this point
    input [31:0] rs1_value_i;
    input [31:0] rs2_value_i;
    
    // Outputs
    output writeback_valid_o;
    output [31:0]  writeback_value_o;


/*
`define FUNCT3_MUL      3'b000
`define FUNCT3_MULH     3'b001
`define FUNCT3_MULHSU   3'b010
`define FUNCT3_MULHU    3'b011
`define FUNCT3_DIV      3'b100
`define FUNCT3_DIVU     3'b101
`define FUNCT3_REM      3'b110
`define FUNCT3_REMU     3'b111*/

endmodule
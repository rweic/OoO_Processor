module core ();

endmodule
/* Core */
module core ();


endmodule